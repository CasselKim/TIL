module main();											
	parameter read_filename = "./proj3-input1.txt";		
	parameter N = 10403;
	parameter e = 71;
	
	wire [6:0] 	 ascii_6783_000,	ascii_6783_001, ascii_6783_002, ascii_6783_003,								
				 ascii_6783_004,	ascii_6783_005,	ascii_6783_006,	ascii_6783_007,				
				 ascii_6783_008,	ascii_6783_009,	ascii_6783_010,	ascii_6783_011,				
				 ascii_6783_012,	ascii_6783_013,	ascii_6783_014,	ascii_6783_015,				
				 ascii_6783_016,	ascii_6783_017,	ascii_6783_018,	ascii_6783_019,				
				 ascii_6783_020,	ascii_6783_021,	ascii_6783_022,	ascii_6783_023,				
				 ascii_6783_024,	ascii_6783_025,	ascii_6783_026,	ascii_6783_027,				
				 ascii_6783_028,	ascii_6783_029,	ascii_6783_030,	ascii_6783_031,				
				 ascii_6783_032,	ascii_6783_033,	ascii_6783_034,	ascii_6783_035,				
				 ascii_6783_036,	ascii_6783_037,	ascii_6783_038,	ascii_6783_039,				
				 ascii_6783_040,	ascii_6783_041,	ascii_6783_042,	ascii_6783_043,				
				 ascii_6783_044,	ascii_6783_045,	ascii_6783_046,	ascii_6783_047,				
				 ascii_6783_048,	ascii_6783_049,	ascii_6783_050,	ascii_6783_051,				
				 ascii_6783_052,	ascii_6783_053,	ascii_6783_054,	ascii_6783_055,				
				 ascii_6783_056,	ascii_6783_057,	ascii_6783_058,	ascii_6783_059,				
				 ascii_6783_060,	ascii_6783_061,	ascii_6783_062,	ascii_6783_063,				
				 ascii_6783_064,	ascii_6783_065,	ascii_6783_066,	ascii_6783_067,				
				 ascii_6783_068,	ascii_6783_069,	ascii_6783_070,	ascii_6783_071,				
				 ascii_6783_072,	ascii_6783_073,	ascii_6783_074,	ascii_6783_075,				
				 ascii_6783_076,	ascii_6783_077,	ascii_6783_078,	ascii_6783_079,				
				 ascii_6783_080,	ascii_6783_081,	ascii_6783_082,	ascii_6783_083,				
				 ascii_6783_084,	ascii_6783_085,	ascii_6783_086,	ascii_6783_087,				
				 ascii_6783_088,	ascii_6783_089,	ascii_6783_090,	ascii_6783_091,				
				 ascii_6783_092,	ascii_6783_093,	ascii_6783_094,	ascii_6783_095,				
				 ascii_6783_096,	ascii_6783_097,	ascii_6783_098,	ascii_6783_099,				
				 ascii_6783_100,	ascii_6783_101,	ascii_6783_102,	ascii_6783_103,				
				 ascii_6783_104,	ascii_6783_105,	ascii_6783_106,	ascii_6783_107,				
				 ascii_6783_108,	ascii_6783_109,	ascii_6783_110,	ascii_6783_111,				
				 ascii_6783_112,	ascii_6783_113,	ascii_6783_114,	ascii_6783_115,				
				 ascii_6783_116,	ascii_6783_117,	ascii_6783_118,	ascii_6783_119,				
				 ascii_6783_120,	ascii_6783_121,	ascii_6783_122,	ascii_6783_123,				
				 ascii_6783_124,	ascii_6783_125,	ascii_6783_126,	ascii_6783_127,				
				 ascii_6783_128,	ascii_6783_129,	ascii_6783_130,	ascii_6783_131,				
				 ascii_6783_132,	ascii_6783_133,	ascii_6783_134,	ascii_6783_135,				
				 ascii_6783_136,	ascii_6783_137,	ascii_6783_138,	ascii_6783_139,				
				 ascii_6783_140,	ascii_6783_141,	ascii_6783_142,	ascii_6783_143,				
				 ascii_6783_144,	ascii_6783_145;
	wire [5:0]   tgBASE_6783_000,	tgBASE_6783_001,    tgBASE_6783_002,    tgBASE_6783_003,							
				 tgBASE_6783_004,	tgBASE_6783_005,	tgBASE_6783_006,	tgBASE_6783_007,	
				 tgBASE_6783_008,	tgBASE_6783_009,	tgBASE_6783_010,	tgBASE_6783_011,	
				 tgBASE_6783_012,	tgBASE_6783_013,	tgBASE_6783_014,	tgBASE_6783_015,	
				 tgBASE_6783_016,	tgBASE_6783_017,	tgBASE_6783_018,	tgBASE_6783_019,	
				 tgBASE_6783_020,	tgBASE_6783_021,	tgBASE_6783_022,	tgBASE_6783_023,	
				 tgBASE_6783_024,	tgBASE_6783_025,	tgBASE_6783_026,	tgBASE_6783_027,	
				 tgBASE_6783_028,	tgBASE_6783_029,	tgBASE_6783_030,	tgBASE_6783_031,	
				 tgBASE_6783_032,	tgBASE_6783_033,	tgBASE_6783_034,	tgBASE_6783_035,	
				 tgBASE_6783_036,	tgBASE_6783_037,	tgBASE_6783_038,	tgBASE_6783_039,	
				 tgBASE_6783_040,	tgBASE_6783_041,	tgBASE_6783_042,	tgBASE_6783_043,	
				 tgBASE_6783_044,	tgBASE_6783_045,	tgBASE_6783_046,	tgBASE_6783_047,	
				 tgBASE_6783_048,	tgBASE_6783_049,	tgBASE_6783_050,	tgBASE_6783_051,	
				 tgBASE_6783_052,	tgBASE_6783_053,	tgBASE_6783_054,	tgBASE_6783_055,	
				 tgBASE_6783_056,	tgBASE_6783_057,	tgBASE_6783_058,	tgBASE_6783_059,	
				 tgBASE_6783_060,	tgBASE_6783_061,	tgBASE_6783_062,	tgBASE_6783_063,	
				 tgBASE_6783_064,	tgBASE_6783_065,	tgBASE_6783_066,	tgBASE_6783_067,	
				 tgBASE_6783_068,	tgBASE_6783_069,	tgBASE_6783_070,	tgBASE_6783_071,	
				 tgBASE_6783_072,	tgBASE_6783_073,	tgBASE_6783_074,	tgBASE_6783_075,	
				 tgBASE_6783_076,	tgBASE_6783_077,	tgBASE_6783_078,	tgBASE_6783_079,	
				 tgBASE_6783_080,	tgBASE_6783_081,	tgBASE_6783_082,	tgBASE_6783_083,	
				 tgBASE_6783_084,	tgBASE_6783_085,	tgBASE_6783_086,	tgBASE_6783_087,	
				 tgBASE_6783_088,	tgBASE_6783_089,	tgBASE_6783_090,	tgBASE_6783_091,	
				 tgBASE_6783_092,	tgBASE_6783_093,	tgBASE_6783_094,	tgBASE_6783_095,	
				 tgBASE_6783_096,	tgBASE_6783_097,	tgBASE_6783_098,	tgBASE_6783_099,	
				 tgBASE_6783_100,	tgBASE_6783_101,	tgBASE_6783_102,	tgBASE_6783_103,	
				 tgBASE_6783_104,	tgBASE_6783_105,	tgBASE_6783_106,	tgBASE_6783_107,	
				 tgBASE_6783_108,	tgBASE_6783_109,	tgBASE_6783_110,	tgBASE_6783_111,	
				 tgBASE_6783_112,	tgBASE_6783_113,	tgBASE_6783_114,	tgBASE_6783_115,	
				 tgBASE_6783_116,	tgBASE_6783_117,	tgBASE_6783_118,	tgBASE_6783_119,	
				 tgBASE_6783_120,	tgBASE_6783_121,	tgBASE_6783_122,	tgBASE_6783_123,	
				 tgBASE_6783_124,	tgBASE_6783_125,	tgBASE_6783_126,	tgBASE_6783_127,	
				 tgBASE_6783_128,	tgBASE_6783_129,	tgBASE_6783_130,	tgBASE_6783_131,	
				 tgBASE_6783_132,	tgBASE_6783_133,	tgBASE_6783_134,	tgBASE_6783_135,	
				 tgBASE_6783_136,	tgBASE_6783_137,	tgBASE_6783_138,	tgBASE_6783_139,	
				 tgBASE_6783_140,	tgBASE_6783_141,	tgBASE_6783_142,	tgBASE_6783_143,	
				 tgBASE_6783_144,	tgBASE_6783_145;
	wire [13:0]  oneBig_6783_000,	oneBig_6783_001,    oneBig_6783_002,    oneBig_6783_003,							
				 oneBig_6783_004,	oneBig_6783_005,	oneBig_6783_006,	oneBig_6783_007,	
				 oneBig_6783_008,	oneBig_6783_009,	oneBig_6783_010,	oneBig_6783_011,	
				 oneBig_6783_012,	oneBig_6783_013,	oneBig_6783_014,	oneBig_6783_015,	
				 oneBig_6783_016,	oneBig_6783_017,	oneBig_6783_018,	oneBig_6783_019,	
				 oneBig_6783_020,	oneBig_6783_021,	oneBig_6783_022,	oneBig_6783_023,	
				 oneBig_6783_024,	oneBig_6783_025,	oneBig_6783_026,	oneBig_6783_027,	
				 oneBig_6783_028,	oneBig_6783_029,	oneBig_6783_030,	oneBig_6783_031,	
				 oneBig_6783_032,	oneBig_6783_033,	oneBig_6783_034,	oneBig_6783_035,	
				 oneBig_6783_036,	oneBig_6783_037,	oneBig_6783_038,	oneBig_6783_039,	
				 oneBig_6783_040,	oneBig_6783_041,	oneBig_6783_042,	oneBig_6783_043,	
				 oneBig_6783_044,	oneBig_6783_045,	oneBig_6783_046,	oneBig_6783_047,	
				 oneBig_6783_048,	oneBig_6783_049,	oneBig_6783_050,	oneBig_6783_051,	
				 oneBig_6783_052,	oneBig_6783_053,	oneBig_6783_054,	oneBig_6783_055,	
				 oneBig_6783_056,	oneBig_6783_057,	oneBig_6783_058,	oneBig_6783_059,	
				 oneBig_6783_060,	oneBig_6783_061,	oneBig_6783_062,	oneBig_6783_063,	
				 oneBig_6783_064,	oneBig_6783_065,	oneBig_6783_066,	oneBig_6783_067,	
				 oneBig_6783_068,	oneBig_6783_069,	oneBig_6783_070,	oneBig_6783_071,	
				 oneBig_6783_072,
				 encrypt_6783_000,	encrypt_6783_001,   encrypt_6783_002,   encrypt_6783_003,							
				 encrypt_6783_004,	encrypt_6783_005,	encrypt_6783_006,	encrypt_6783_007,	
				 encrypt_6783_008,	encrypt_6783_009,	encrypt_6783_010,	encrypt_6783_011,	
				 encrypt_6783_012,	encrypt_6783_013,	encrypt_6783_014,	encrypt_6783_015,	
				 encrypt_6783_016,	encrypt_6783_017,	encrypt_6783_018,	encrypt_6783_019,	
				 encrypt_6783_020,	encrypt_6783_021,	encrypt_6783_022,	encrypt_6783_023,	
				 encrypt_6783_024,	encrypt_6783_025,	encrypt_6783_026,	encrypt_6783_027,	
				 encrypt_6783_028,	encrypt_6783_029,	encrypt_6783_030,	encrypt_6783_031,	
				 encrypt_6783_032,	encrypt_6783_033,	encrypt_6783_034,	encrypt_6783_035,	
				 encrypt_6783_036,	encrypt_6783_037,	encrypt_6783_038,	encrypt_6783_039,	
				 encrypt_6783_040,	encrypt_6783_041,	encrypt_6783_042,	encrypt_6783_043,	
				 encrypt_6783_044,	encrypt_6783_045,	encrypt_6783_046,	encrypt_6783_047,	
				 encrypt_6783_048,	encrypt_6783_049,	encrypt_6783_050,	encrypt_6783_051,	
				 encrypt_6783_052,	encrypt_6783_053,	encrypt_6783_054,	encrypt_6783_055,	
				 encrypt_6783_056,	encrypt_6783_057,	encrypt_6783_058,	encrypt_6783_059,	
				 encrypt_6783_060,	encrypt_6783_061,	encrypt_6783_062,	encrypt_6783_063,	
				 encrypt_6783_064,	encrypt_6783_065,	encrypt_6783_066,	encrypt_6783_067,	
				 encrypt_6783_068,	encrypt_6783_069,	encrypt_6783_070,	encrypt_6783_071,	
				 encrypt_6783_072,
				 DoneBig_6783_000,	DoneBig_6783_001,   DoneBig_6783_002,   DoneBig_6783_003,							
				 DoneBig_6783_004,	DoneBig_6783_005,	DoneBig_6783_006,	DoneBig_6783_007,	
				 DoneBig_6783_008,	DoneBig_6783_009,	DoneBig_6783_010,	DoneBig_6783_011,	
				 DoneBig_6783_012,	DoneBig_6783_013,	DoneBig_6783_014,	DoneBig_6783_015,	
				 DoneBig_6783_016,	DoneBig_6783_017,	DoneBig_6783_018,	DoneBig_6783_019,	
				 DoneBig_6783_020,	DoneBig_6783_021,	DoneBig_6783_022,	DoneBig_6783_023,	
				 DoneBig_6783_024,	DoneBig_6783_025,	DoneBig_6783_026,	DoneBig_6783_027,	
				 DoneBig_6783_028,	DoneBig_6783_029,	DoneBig_6783_030,	DoneBig_6783_031,	
				 DoneBig_6783_032,	DoneBig_6783_033,	DoneBig_6783_034,	DoneBig_6783_035,	
				 DoneBig_6783_036,	DoneBig_6783_037,	DoneBig_6783_038,	DoneBig_6783_039,	
				 DoneBig_6783_040,	DoneBig_6783_041,	DoneBig_6783_042,	DoneBig_6783_043,	
				 DoneBig_6783_044,	DoneBig_6783_045,	DoneBig_6783_046,	DoneBig_6783_047,	
				 DoneBig_6783_048,	DoneBig_6783_049,	DoneBig_6783_050,	DoneBig_6783_051,	
				 DoneBig_6783_052,	DoneBig_6783_053,	DoneBig_6783_054,	DoneBig_6783_055,	
				 DoneBig_6783_056,	DoneBig_6783_057,	DoneBig_6783_058,	DoneBig_6783_059,	
				 DoneBig_6783_060,	DoneBig_6783_061,	DoneBig_6783_062,	DoneBig_6783_063,	
				 DoneBig_6783_064,	DoneBig_6783_065,	DoneBig_6783_066,	DoneBig_6783_067,	
				 DoneBig_6783_068,	DoneBig_6783_069,	DoneBig_6783_070,	DoneBig_6783_071,	
				 DoneBig_6783_072;				

				

	reg [1022:0] ascii_IN;										
	integer fp;										
											
	ascii_IN_to_ascii_6783_ u1(ascii_IN, 										
				 ascii_6783_000,	ascii_6783_001, ascii_6783_002, ascii_6783_003,						
				 ascii_6783_004,	ascii_6783_005,	ascii_6783_006,	ascii_6783_007,				
				 ascii_6783_008,	ascii_6783_009,	ascii_6783_010,	ascii_6783_011,				
				 ascii_6783_012,	ascii_6783_013,	ascii_6783_014,	ascii_6783_015,				
				 ascii_6783_016,	ascii_6783_017,	ascii_6783_018,	ascii_6783_019,				
				 ascii_6783_020,	ascii_6783_021,	ascii_6783_022,	ascii_6783_023,				
				 ascii_6783_024,	ascii_6783_025,	ascii_6783_026,	ascii_6783_027,				
				 ascii_6783_028,	ascii_6783_029,	ascii_6783_030,	ascii_6783_031,				
				 ascii_6783_032,	ascii_6783_033,	ascii_6783_034,	ascii_6783_035,				
				 ascii_6783_036,	ascii_6783_037,	ascii_6783_038,	ascii_6783_039,				
				 ascii_6783_040,	ascii_6783_041,	ascii_6783_042,	ascii_6783_043,				
				 ascii_6783_044,	ascii_6783_045,	ascii_6783_046,	ascii_6783_047,				
				 ascii_6783_048,	ascii_6783_049,	ascii_6783_050,	ascii_6783_051,				
				 ascii_6783_052,	ascii_6783_053,	ascii_6783_054,	ascii_6783_055,				
				 ascii_6783_056,	ascii_6783_057,	ascii_6783_058,	ascii_6783_059,				
				 ascii_6783_060,	ascii_6783_061,	ascii_6783_062,	ascii_6783_063,				
				 ascii_6783_064,	ascii_6783_065,	ascii_6783_066,	ascii_6783_067,				
				 ascii_6783_068,	ascii_6783_069,	ascii_6783_070,	ascii_6783_071,				
				 ascii_6783_072,	ascii_6783_073,	ascii_6783_074,	ascii_6783_075,				
				 ascii_6783_076,	ascii_6783_077,	ascii_6783_078,	ascii_6783_079,				
				 ascii_6783_080,	ascii_6783_081,	ascii_6783_082,	ascii_6783_083,				
				 ascii_6783_084,	ascii_6783_085,	ascii_6783_086,	ascii_6783_087,				
				 ascii_6783_088,	ascii_6783_089,	ascii_6783_090,	ascii_6783_091,				
				 ascii_6783_092,	ascii_6783_093,	ascii_6783_094,	ascii_6783_095,				
				 ascii_6783_096,	ascii_6783_097,	ascii_6783_098,	ascii_6783_099,				
				 ascii_6783_100,	ascii_6783_101,	ascii_6783_102,	ascii_6783_103,				
				 ascii_6783_104,	ascii_6783_105,	ascii_6783_106,	ascii_6783_107,				
				 ascii_6783_108,	ascii_6783_109,	ascii_6783_110,	ascii_6783_111,				
				 ascii_6783_112,	ascii_6783_113,	ascii_6783_114,	ascii_6783_115,				
				 ascii_6783_116,	ascii_6783_117,	ascii_6783_118,	ascii_6783_119,				
				 ascii_6783_120,	ascii_6783_121,	ascii_6783_122,	ascii_6783_123,				
				 ascii_6783_124,	ascii_6783_125,	ascii_6783_126,	ascii_6783_127,				
				 ascii_6783_128,	ascii_6783_129,	ascii_6783_130,	ascii_6783_131,				
				 ascii_6783_132,	ascii_6783_133,	ascii_6783_134,	ascii_6783_135,				
				 ascii_6783_136,	ascii_6783_137,	ascii_6783_138,	ascii_6783_139,				
				 ascii_6783_140,	ascii_6783_141,	ascii_6783_142,	ascii_6783_143,				
				 ascii_6783_144,	ascii_6783_145);						
											
	ascii7b_to_tgbase64 u2(
				 ascii_6783_000,	ascii_6783_001, ascii_6783_002, ascii_6783_003,									
				 ascii_6783_004,	ascii_6783_005,	ascii_6783_006,	ascii_6783_007,				
				 ascii_6783_008,	ascii_6783_009,	ascii_6783_010,	ascii_6783_011,				
				 ascii_6783_012,	ascii_6783_013,	ascii_6783_014,	ascii_6783_015,				
				 ascii_6783_016,	ascii_6783_017,	ascii_6783_018,	ascii_6783_019,				
				 ascii_6783_020,	ascii_6783_021,	ascii_6783_022,	ascii_6783_023,				
				 ascii_6783_024,	ascii_6783_025,	ascii_6783_026,	ascii_6783_027,				
				 ascii_6783_028,	ascii_6783_029,	ascii_6783_030,	ascii_6783_031,				
				 ascii_6783_032,	ascii_6783_033,	ascii_6783_034,	ascii_6783_035,				
				 ascii_6783_036,	ascii_6783_037,	ascii_6783_038,	ascii_6783_039,				
				 ascii_6783_040,	ascii_6783_041,	ascii_6783_042,	ascii_6783_043,				
				 ascii_6783_044,	ascii_6783_045,	ascii_6783_046,	ascii_6783_047,				
				 ascii_6783_048,	ascii_6783_049,	ascii_6783_050,	ascii_6783_051,				
				 ascii_6783_052,	ascii_6783_053,	ascii_6783_054,	ascii_6783_055,				
				 ascii_6783_056,	ascii_6783_057,	ascii_6783_058,	ascii_6783_059,				
				 ascii_6783_060,	ascii_6783_061,	ascii_6783_062,	ascii_6783_063,				
				 ascii_6783_064,	ascii_6783_065,	ascii_6783_066,	ascii_6783_067,				
				 ascii_6783_068,	ascii_6783_069,	ascii_6783_070,	ascii_6783_071,				
				 ascii_6783_072,	ascii_6783_073,	ascii_6783_074,	ascii_6783_075,				
				 ascii_6783_076,	ascii_6783_077,	ascii_6783_078,	ascii_6783_079,				
				 ascii_6783_080,	ascii_6783_081,	ascii_6783_082,	ascii_6783_083,				
				 ascii_6783_084,	ascii_6783_085,	ascii_6783_086,	ascii_6783_087,				
				 ascii_6783_088,	ascii_6783_089,	ascii_6783_090,	ascii_6783_091,				
				 ascii_6783_092,	ascii_6783_093,	ascii_6783_094,	ascii_6783_095,				
				 ascii_6783_096,	ascii_6783_097,	ascii_6783_098,	ascii_6783_099,				
				 ascii_6783_100,	ascii_6783_101,	ascii_6783_102,	ascii_6783_103,				
				 ascii_6783_104,	ascii_6783_105,	ascii_6783_106,	ascii_6783_107,				
				 ascii_6783_108,	ascii_6783_109,	ascii_6783_110,	ascii_6783_111,				
				 ascii_6783_112,	ascii_6783_113,	ascii_6783_114,	ascii_6783_115,				
				 ascii_6783_116,	ascii_6783_117,	ascii_6783_118,	ascii_6783_119,				
				 ascii_6783_120,	ascii_6783_121,	ascii_6783_122,	ascii_6783_123,				
				 ascii_6783_124,	ascii_6783_125,	ascii_6783_126,	ascii_6783_127,				
				 ascii_6783_128,	ascii_6783_129,	ascii_6783_130,	ascii_6783_131,				
				 ascii_6783_132,	ascii_6783_133,	ascii_6783_134,	ascii_6783_135,				
				 ascii_6783_136,	ascii_6783_137,	ascii_6783_138,	ascii_6783_139,				
				 ascii_6783_140,	ascii_6783_141,	ascii_6783_142,	ascii_6783_143,				
				 ascii_6783_144,	ascii_6783_145,
				 tgBASE_6783_000,	tgBASE_6783_001,    tgBASE_6783_002,    tgBASE_6783_003,							
				 tgBASE_6783_004,	tgBASE_6783_005,	tgBASE_6783_006,	tgBASE_6783_007,	
				 tgBASE_6783_008,	tgBASE_6783_009,	tgBASE_6783_010,	tgBASE_6783_011,	
				 tgBASE_6783_012,	tgBASE_6783_013,	tgBASE_6783_014,	tgBASE_6783_015,	
				 tgBASE_6783_016,	tgBASE_6783_017,	tgBASE_6783_018,	tgBASE_6783_019,	
				 tgBASE_6783_020,	tgBASE_6783_021,	tgBASE_6783_022,	tgBASE_6783_023,	
				 tgBASE_6783_024,	tgBASE_6783_025,	tgBASE_6783_026,	tgBASE_6783_027,	
				 tgBASE_6783_028,	tgBASE_6783_029,	tgBASE_6783_030,	tgBASE_6783_031,	
				 tgBASE_6783_032,	tgBASE_6783_033,	tgBASE_6783_034,	tgBASE_6783_035,	
				 tgBASE_6783_036,	tgBASE_6783_037,	tgBASE_6783_038,	tgBASE_6783_039,	
				 tgBASE_6783_040,	tgBASE_6783_041,	tgBASE_6783_042,	tgBASE_6783_043,	
				 tgBASE_6783_044,	tgBASE_6783_045,	tgBASE_6783_046,	tgBASE_6783_047,	
				 tgBASE_6783_048,	tgBASE_6783_049,	tgBASE_6783_050,	tgBASE_6783_051,	
				 tgBASE_6783_052,	tgBASE_6783_053,	tgBASE_6783_054,	tgBASE_6783_055,	
				 tgBASE_6783_056,	tgBASE_6783_057,	tgBASE_6783_058,	tgBASE_6783_059,	
				 tgBASE_6783_060,	tgBASE_6783_061,	tgBASE_6783_062,	tgBASE_6783_063,	
				 tgBASE_6783_064,	tgBASE_6783_065,	tgBASE_6783_066,	tgBASE_6783_067,	
				 tgBASE_6783_068,	tgBASE_6783_069,	tgBASE_6783_070,	tgBASE_6783_071,	
				 tgBASE_6783_072,	tgBASE_6783_073,	tgBASE_6783_074,	tgBASE_6783_075,	
				 tgBASE_6783_076,	tgBASE_6783_077,	tgBASE_6783_078,	tgBASE_6783_079,	
				 tgBASE_6783_080,	tgBASE_6783_081,	tgBASE_6783_082,	tgBASE_6783_083,	
				 tgBASE_6783_084,	tgBASE_6783_085,	tgBASE_6783_086,	tgBASE_6783_087,	
				 tgBASE_6783_088,	tgBASE_6783_089,	tgBASE_6783_090,	tgBASE_6783_091,	
				 tgBASE_6783_092,	tgBASE_6783_093,	tgBASE_6783_094,	tgBASE_6783_095,	
				 tgBASE_6783_096,	tgBASE_6783_097,	tgBASE_6783_098,	tgBASE_6783_099,	
				 tgBASE_6783_100,	tgBASE_6783_101,	tgBASE_6783_102,	tgBASE_6783_103,	
				 tgBASE_6783_104,	tgBASE_6783_105,	tgBASE_6783_106,	tgBASE_6783_107,	
				 tgBASE_6783_108,	tgBASE_6783_109,	tgBASE_6783_110,	tgBASE_6783_111,	
				 tgBASE_6783_112,	tgBASE_6783_113,	tgBASE_6783_114,	tgBASE_6783_115,	
				 tgBASE_6783_116,	tgBASE_6783_117,	tgBASE_6783_118,	tgBASE_6783_119,	
				 tgBASE_6783_120,	tgBASE_6783_121,	tgBASE_6783_122,	tgBASE_6783_123,	
				 tgBASE_6783_124,	tgBASE_6783_125,	tgBASE_6783_126,	tgBASE_6783_127,	
				 tgBASE_6783_128,	tgBASE_6783_129,	tgBASE_6783_130,	tgBASE_6783_131,	
				 tgBASE_6783_132,	tgBASE_6783_133,	tgBASE_6783_134,	tgBASE_6783_135,	
				 tgBASE_6783_136,	tgBASE_6783_137,	tgBASE_6783_138,	tgBASE_6783_139,	
				 tgBASE_6783_140,	tgBASE_6783_141,	tgBASE_6783_142,	tgBASE_6783_143,	
				 tgBASE_6783_144,	tgBASE_6783_145);
				 
	two_tgbase_to_one_big_number u3(
				 tgBASE_6783_000,	tgBASE_6783_001,    tgBASE_6783_002,    tgBASE_6783_003,							
				 tgBASE_6783_004,	tgBASE_6783_005,	tgBASE_6783_006,	tgBASE_6783_007,	
				 tgBASE_6783_008,	tgBASE_6783_009,	tgBASE_6783_010,	tgBASE_6783_011,	
				 tgBASE_6783_012,	tgBASE_6783_013,	tgBASE_6783_014,	tgBASE_6783_015,	
				 tgBASE_6783_016,	tgBASE_6783_017,	tgBASE_6783_018,	tgBASE_6783_019,	
				 tgBASE_6783_020,	tgBASE_6783_021,	tgBASE_6783_022,	tgBASE_6783_023,	
				 tgBASE_6783_024,	tgBASE_6783_025,	tgBASE_6783_026,	tgBASE_6783_027,	
				 tgBASE_6783_028,	tgBASE_6783_029,	tgBASE_6783_030,	tgBASE_6783_031,	
				 tgBASE_6783_032,	tgBASE_6783_033,	tgBASE_6783_034,	tgBASE_6783_035,	
				 tgBASE_6783_036,	tgBASE_6783_037,	tgBASE_6783_038,	tgBASE_6783_039,	
				 tgBASE_6783_040,	tgBASE_6783_041,	tgBASE_6783_042,	tgBASE_6783_043,	
				 tgBASE_6783_044,	tgBASE_6783_045,	tgBASE_6783_046,	tgBASE_6783_047,	
				 tgBASE_6783_048,	tgBASE_6783_049,	tgBASE_6783_050,	tgBASE_6783_051,	
				 tgBASE_6783_052,	tgBASE_6783_053,	tgBASE_6783_054,	tgBASE_6783_055,	
				 tgBASE_6783_056,	tgBASE_6783_057,	tgBASE_6783_058,	tgBASE_6783_059,	
				 tgBASE_6783_060,	tgBASE_6783_061,	tgBASE_6783_062,	tgBASE_6783_063,	
				 tgBASE_6783_064,	tgBASE_6783_065,	tgBASE_6783_066,	tgBASE_6783_067,	
				 tgBASE_6783_068,	tgBASE_6783_069,	tgBASE_6783_070,	tgBASE_6783_071,	
				 tgBASE_6783_072,	tgBASE_6783_073,	tgBASE_6783_074,	tgBASE_6783_075,	
				 tgBASE_6783_076,	tgBASE_6783_077,	tgBASE_6783_078,	tgBASE_6783_079,	
				 tgBASE_6783_080,	tgBASE_6783_081,	tgBASE_6783_082,	tgBASE_6783_083,	
				 tgBASE_6783_084,	tgBASE_6783_085,	tgBASE_6783_086,	tgBASE_6783_087,	
				 tgBASE_6783_088,	tgBASE_6783_089,	tgBASE_6783_090,	tgBASE_6783_091,	
				 tgBASE_6783_092,	tgBASE_6783_093,	tgBASE_6783_094,	tgBASE_6783_095,	
				 tgBASE_6783_096,	tgBASE_6783_097,	tgBASE_6783_098,	tgBASE_6783_099,	
				 tgBASE_6783_100,	tgBASE_6783_101,	tgBASE_6783_102,	tgBASE_6783_103,	
				 tgBASE_6783_104,	tgBASE_6783_105,	tgBASE_6783_106,	tgBASE_6783_107,	
				 tgBASE_6783_108,	tgBASE_6783_109,	tgBASE_6783_110,	tgBASE_6783_111,	
				 tgBASE_6783_112,	tgBASE_6783_113,	tgBASE_6783_114,	tgBASE_6783_115,	
				 tgBASE_6783_116,	tgBASE_6783_117,	tgBASE_6783_118,	tgBASE_6783_119,	
				 tgBASE_6783_120,	tgBASE_6783_121,	tgBASE_6783_122,	tgBASE_6783_123,	
				 tgBASE_6783_124,	tgBASE_6783_125,	tgBASE_6783_126,	tgBASE_6783_127,	
				 tgBASE_6783_128,	tgBASE_6783_129,	tgBASE_6783_130,	tgBASE_6783_131,	
				 tgBASE_6783_132,	tgBASE_6783_133,	tgBASE_6783_134,	tgBASE_6783_135,	
				 tgBASE_6783_136,	tgBASE_6783_137,	tgBASE_6783_138,	tgBASE_6783_139,	
				 tgBASE_6783_140,	tgBASE_6783_141,	tgBASE_6783_142,	tgBASE_6783_143,	
				 tgBASE_6783_144,	tgBASE_6783_145,
				 oneBig_6783_000,	oneBig_6783_001,    oneBig_6783_002,    oneBig_6783_003,							
				 oneBig_6783_004,	oneBig_6783_005,	oneBig_6783_006,	oneBig_6783_007,	
				 oneBig_6783_008,	oneBig_6783_009,	oneBig_6783_010,	oneBig_6783_011,	
				 oneBig_6783_012,	oneBig_6783_013,	oneBig_6783_014,	oneBig_6783_015,	
				 oneBig_6783_016,	oneBig_6783_017,	oneBig_6783_018,	oneBig_6783_019,	
				 oneBig_6783_020,	oneBig_6783_021,	oneBig_6783_022,	oneBig_6783_023,	
				 oneBig_6783_024,	oneBig_6783_025,	oneBig_6783_026,	oneBig_6783_027,	
				 oneBig_6783_028,	oneBig_6783_029,	oneBig_6783_030,	oneBig_6783_031,	
				 oneBig_6783_032,	oneBig_6783_033,	oneBig_6783_034,	oneBig_6783_035,	
				 oneBig_6783_036,	oneBig_6783_037,	oneBig_6783_038,	oneBig_6783_039,	
				 oneBig_6783_040,	oneBig_6783_041,	oneBig_6783_042,	oneBig_6783_043,	
				 oneBig_6783_044,	oneBig_6783_045,	oneBig_6783_046,	oneBig_6783_047,	
				 oneBig_6783_048,	oneBig_6783_049,	oneBig_6783_050,	oneBig_6783_051,	
				 oneBig_6783_052,	oneBig_6783_053,	oneBig_6783_054,	oneBig_6783_055,	
				 oneBig_6783_056,	oneBig_6783_057,	oneBig_6783_058,	oneBig_6783_059,	
				 oneBig_6783_060,	oneBig_6783_061,	oneBig_6783_062,	oneBig_6783_063,	
				 oneBig_6783_064,	oneBig_6783_065,	oneBig_6783_066,	oneBig_6783_067,	
				 oneBig_6783_068,	oneBig_6783_069,	oneBig_6783_070,	oneBig_6783_071,	
				 oneBig_6783_072);
	
	rsa_encryption u4(N, e,
				 oneBig_6783_000,	oneBig_6783_001,    oneBig_6783_002,    oneBig_6783_003,							
				 oneBig_6783_004,	oneBig_6783_005,	oneBig_6783_006,	oneBig_6783_007,	
				 oneBig_6783_008,	oneBig_6783_009,	oneBig_6783_010,	oneBig_6783_011,	
				 oneBig_6783_012,	oneBig_6783_013,	oneBig_6783_014,	oneBig_6783_015,	
				 oneBig_6783_016,	oneBig_6783_017,	oneBig_6783_018,	oneBig_6783_019,	
				 oneBig_6783_020,	oneBig_6783_021,	oneBig_6783_022,	oneBig_6783_023,	
				 oneBig_6783_024,	oneBig_6783_025,	oneBig_6783_026,	oneBig_6783_027,	
				 oneBig_6783_028,	oneBig_6783_029,	oneBig_6783_030,	oneBig_6783_031,	
				 oneBig_6783_032,	oneBig_6783_033,	oneBig_6783_034,	oneBig_6783_035,	
				 oneBig_6783_036,	oneBig_6783_037,	oneBig_6783_038,	oneBig_6783_039,	
				 oneBig_6783_040,	oneBig_6783_041,	oneBig_6783_042,	oneBig_6783_043,	
				 oneBig_6783_044,	oneBig_6783_045,	oneBig_6783_046,	oneBig_6783_047,	
				 oneBig_6783_048,	oneBig_6783_049,	oneBig_6783_050,	oneBig_6783_051,	
				 oneBig_6783_052,	oneBig_6783_053,	oneBig_6783_054,	oneBig_6783_055,	
				 oneBig_6783_056,	oneBig_6783_057,	oneBig_6783_058,	oneBig_6783_059,	
				 oneBig_6783_060,	oneBig_6783_061,	oneBig_6783_062,	oneBig_6783_063,	
				 oneBig_6783_064,	oneBig_6783_065,	oneBig_6783_066,	oneBig_6783_067,	
				 oneBig_6783_068,	oneBig_6783_069,	oneBig_6783_070,	oneBig_6783_071,	
				 oneBig_6783_072,
				 encrypt_6783_000,	encrypt_6783_001,   encrypt_6783_002,   encrypt_6783_003,							
				 encrypt_6783_004,	encrypt_6783_005,	encrypt_6783_006,	encrypt_6783_007,	
				 encrypt_6783_008,	encrypt_6783_009,	encrypt_6783_010,	encrypt_6783_011,	
				 encrypt_6783_012,	encrypt_6783_013,	encrypt_6783_014,	encrypt_6783_015,	
				 encrypt_6783_016,	encrypt_6783_017,	encrypt_6783_018,	encrypt_6783_019,	
				 encrypt_6783_020,	encrypt_6783_021,	encrypt_6783_022,	encrypt_6783_023,	
				 encrypt_6783_024,	encrypt_6783_025,	encrypt_6783_026,	encrypt_6783_027,	
				 encrypt_6783_028,	encrypt_6783_029,	encrypt_6783_030,	encrypt_6783_031,	
				 encrypt_6783_032,	encrypt_6783_033,	encrypt_6783_034,	encrypt_6783_035,	
				 encrypt_6783_036,	encrypt_6783_037,	encrypt_6783_038,	encrypt_6783_039,	
				 encrypt_6783_040,	encrypt_6783_041,	encrypt_6783_042,	encrypt_6783_043,	
				 encrypt_6783_044,	encrypt_6783_045,	encrypt_6783_046,	encrypt_6783_047,	
				 encrypt_6783_048,	encrypt_6783_049,	encrypt_6783_050,	encrypt_6783_051,	
				 encrypt_6783_052,	encrypt_6783_053,	encrypt_6783_054,	encrypt_6783_055,	
				 encrypt_6783_056,	encrypt_6783_057,	encrypt_6783_058,	encrypt_6783_059,	
				 encrypt_6783_060,	encrypt_6783_061,	encrypt_6783_062,	encrypt_6783_063,	
				 encrypt_6783_064,	encrypt_6783_065,	encrypt_6783_066,	encrypt_6783_067,	
				 encrypt_6783_068,	encrypt_6783_069,	encrypt_6783_070,	encrypt_6783_071,	
				 encrypt_6783_072);
				 
	rsa_decryption u5(N,e,
				 encrypt_6783_000,	encrypt_6783_001,   encrypt_6783_002,   encrypt_6783_003,							
				 encrypt_6783_004,	encrypt_6783_005,	encrypt_6783_006,	encrypt_6783_007,	
				 encrypt_6783_008,	encrypt_6783_009,	encrypt_6783_010,	encrypt_6783_011,	
				 encrypt_6783_012,	encrypt_6783_013,	encrypt_6783_014,	encrypt_6783_015,	
				 encrypt_6783_016,	encrypt_6783_017,	encrypt_6783_018,	encrypt_6783_019,	
				 encrypt_6783_020,	encrypt_6783_021,	encrypt_6783_022,	encrypt_6783_023,	
				 encrypt_6783_024,	encrypt_6783_025,	encrypt_6783_026,	encrypt_6783_027,	
				 encrypt_6783_028,	encrypt_6783_029,	encrypt_6783_030,	encrypt_6783_031,	
				 encrypt_6783_032,	encrypt_6783_033,	encrypt_6783_034,	encrypt_6783_035,	
				 encrypt_6783_036,	encrypt_6783_037,	encrypt_6783_038,	encrypt_6783_039,	
				 encrypt_6783_040,	encrypt_6783_041,	encrypt_6783_042,	encrypt_6783_043,	
				 encrypt_6783_044,	encrypt_6783_045,	encrypt_6783_046,	encrypt_6783_047,	
				 encrypt_6783_048,	encrypt_6783_049,	encrypt_6783_050,	encrypt_6783_051,	
				 encrypt_6783_052,	encrypt_6783_053,	encrypt_6783_054,	encrypt_6783_055,	
				 encrypt_6783_056,	encrypt_6783_057,	encrypt_6783_058,	encrypt_6783_059,	
				 encrypt_6783_060,	encrypt_6783_061,	encrypt_6783_062,	encrypt_6783_063,	
				 encrypt_6783_064,	encrypt_6783_065,	encrypt_6783_066,	encrypt_6783_067,	
				 encrypt_6783_068,	encrypt_6783_069,	encrypt_6783_070,	encrypt_6783_071,	
				 encrypt_6783_072,
				 DoneBig_6783_000,	DoneBig_6783_001,   DoneBig_6783_002,   DoneBig_6783_003,							
				 DoneBig_6783_004,	DoneBig_6783_005,	DoneBig_6783_006,	DoneBig_6783_007,	
				 DoneBig_6783_008,	DoneBig_6783_009,	DoneBig_6783_010,	DoneBig_6783_011,	
				 DoneBig_6783_012,	DoneBig_6783_013,	DoneBig_6783_014,	DoneBig_6783_015,	
				 DoneBig_6783_016,	DoneBig_6783_017,	DoneBig_6783_018,	DoneBig_6783_019,	
				 DoneBig_6783_020,	DoneBig_6783_021,	DoneBig_6783_022,	DoneBig_6783_023,	
				 DoneBig_6783_024,	DoneBig_6783_025,	DoneBig_6783_026,	DoneBig_6783_027,	
				 DoneBig_6783_028,	DoneBig_6783_029,	DoneBig_6783_030,	DoneBig_6783_031,	
				 DoneBig_6783_032,	DoneBig_6783_033,	DoneBig_6783_034,	DoneBig_6783_035,	
				 DoneBig_6783_036,	DoneBig_6783_037,	DoneBig_6783_038,	DoneBig_6783_039,	
				 DoneBig_6783_040,	DoneBig_6783_041,	DoneBig_6783_042,	DoneBig_6783_043,	
				 DoneBig_6783_044,	DoneBig_6783_045,	DoneBig_6783_046,	DoneBig_6783_047,	
				 DoneBig_6783_048,	DoneBig_6783_049,	DoneBig_6783_050,	DoneBig_6783_051,	
				 DoneBig_6783_052,	DoneBig_6783_053,	DoneBig_6783_054,	DoneBig_6783_055,	
				 DoneBig_6783_056,	DoneBig_6783_057,	DoneBig_6783_058,	DoneBig_6783_059,	
				 DoneBig_6783_060,	DoneBig_6783_061,	DoneBig_6783_062,	DoneBig_6783_063,	
				 DoneBig_6783_064,	DoneBig_6783_065,	DoneBig_6783_066,	DoneBig_6783_067,	
				 DoneBig_6783_068,	DoneBig_6783_069,	DoneBig_6783_070,	DoneBig_6783_071,	
				 DoneBig_6783_072);				

	
	initial begin										
		fp = $fopen(read_filename, "r");									
		if(!fp) begin									
			$display("read Binary : Open error!\n");								
			$finish;								
		end									
		
		$display("input file : %s\n", read_filename);									
		$fscanf(fp,"%b",ascii_IN);									
		$fclose(fp);									
	end										
	
endmodule											