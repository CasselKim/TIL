module ascii_IN_to_ascii_6783_(								
	input [1022:0] ascii_IN,							
	output [6:0] ascii_6783_000,	ascii_6783_001,  ascii_6783_002,  ascii_6783_003,						
				 ascii_6783_004,	ascii_6783_005,	ascii_6783_006,	ascii_6783_007,	
				 ascii_6783_008,	ascii_6783_009,	ascii_6783_010,	ascii_6783_011,	
				 ascii_6783_012,	ascii_6783_013,	ascii_6783_014,	ascii_6783_015,	
				 ascii_6783_016,	ascii_6783_017,	ascii_6783_018,	ascii_6783_019,	
				 ascii_6783_020,	ascii_6783_021,	ascii_6783_022,	ascii_6783_023,	
				 ascii_6783_024,	ascii_6783_025,	ascii_6783_026,	ascii_6783_027,	
				 ascii_6783_028,	ascii_6783_029,	ascii_6783_030,	ascii_6783_031,	
				 ascii_6783_032,	ascii_6783_033,	ascii_6783_034,	ascii_6783_035,	
				 ascii_6783_036,	ascii_6783_037,	ascii_6783_038,	ascii_6783_039,	
				 ascii_6783_040,	ascii_6783_041,	ascii_6783_042,	ascii_6783_043,	
				 ascii_6783_044,	ascii_6783_045,	ascii_6783_046,	ascii_6783_047,	
				 ascii_6783_048,	ascii_6783_049,	ascii_6783_050,	ascii_6783_051,	
				 ascii_6783_052,	ascii_6783_053,	ascii_6783_054,	ascii_6783_055,	
				 ascii_6783_056,	ascii_6783_057,	ascii_6783_058,	ascii_6783_059,	
				 ascii_6783_060,	ascii_6783_061,	ascii_6783_062,	ascii_6783_063,	
				 ascii_6783_064,	ascii_6783_065,	ascii_6783_066,	ascii_6783_067,	
				 ascii_6783_068,	ascii_6783_069,	ascii_6783_070,	ascii_6783_071,	
				 ascii_6783_072,	ascii_6783_073,	ascii_6783_074,	ascii_6783_075,	
				 ascii_6783_076,	ascii_6783_077,	ascii_6783_078,	ascii_6783_079,	
				 ascii_6783_080,	ascii_6783_081,	ascii_6783_082,	ascii_6783_083,	
				 ascii_6783_084,	ascii_6783_085,	ascii_6783_086,	ascii_6783_087,	
				 ascii_6783_088,	ascii_6783_089,	ascii_6783_090,	ascii_6783_091,	
				 ascii_6783_092,	ascii_6783_093,	ascii_6783_094,	ascii_6783_095,	
				 ascii_6783_096,	ascii_6783_097,	ascii_6783_098,	ascii_6783_099,	
				 ascii_6783_100,	ascii_6783_101,	ascii_6783_102,	ascii_6783_103,	
				 ascii_6783_104,	ascii_6783_105,	ascii_6783_106,	ascii_6783_107,	
				 ascii_6783_108,	ascii_6783_109,	ascii_6783_110,	ascii_6783_111,	
				 ascii_6783_112,	ascii_6783_113,	ascii_6783_114,	ascii_6783_115,	
				 ascii_6783_116,	ascii_6783_117,	ascii_6783_118,	ascii_6783_119,	
				 ascii_6783_120,	ascii_6783_121,	ascii_6783_122,	ascii_6783_123,	
				 ascii_6783_124,	ascii_6783_125,	ascii_6783_126,	ascii_6783_127,	
				 ascii_6783_128,	ascii_6783_129,	ascii_6783_130,	ascii_6783_131,	
				 ascii_6783_132,	ascii_6783_133,	ascii_6783_134,	ascii_6783_135,	
				 ascii_6783_136,	ascii_6783_137,	ascii_6783_138,	ascii_6783_139,	
				 ascii_6783_140,	ascii_6783_141,	ascii_6783_142,	ascii_6783_143,	
				 ascii_6783_144,	ascii_6783_145			
	);							
								
	integer i;							
	assign ascii_6783_000 =ascii_IN[6:0];							
	assign ascii_6783_001 =ascii_IN[13:7];							
	assign ascii_6783_002 =ascii_IN[20:14];							
	assign ascii_6783_003 =ascii_IN[27:21];							
	assign ascii_6783_004 =ascii_IN[34:28];							
	assign ascii_6783_005 =ascii_IN[41:35];							
	assign ascii_6783_006 =ascii_IN[48:42];							
	assign ascii_6783_007 =ascii_IN[55:49];							
	assign ascii_6783_008 =ascii_IN[62:56];							
	assign ascii_6783_009 =ascii_IN[69:63];							
	assign ascii_6783_010 =ascii_IN[76:70];							
	assign ascii_6783_011 =ascii_IN[83:77];							
	assign ascii_6783_012 =ascii_IN[90:84];							
	assign ascii_6783_013 =ascii_IN[97:91];							
	assign ascii_6783_014 =ascii_IN[104:98];							
	assign ascii_6783_015 =ascii_IN[111:105];							
	assign ascii_6783_016 =ascii_IN[118:112];							
	assign ascii_6783_017 =ascii_IN[125:119];							
	assign ascii_6783_018 =ascii_IN[132:126];							
	assign ascii_6783_019 =ascii_IN[139:133];							
	assign ascii_6783_020 =ascii_IN[146:140];							
	assign ascii_6783_021 =ascii_IN[153:147];							
	assign ascii_6783_022 =ascii_IN[160:154];							
	assign ascii_6783_023 =ascii_IN[167:161];							
	assign ascii_6783_024 =ascii_IN[174:168];							
	assign ascii_6783_025 =ascii_IN[181:175];							
	assign ascii_6783_026 =ascii_IN[188:182];							
	assign ascii_6783_027 =ascii_IN[195:189];							
	assign ascii_6783_028 =ascii_IN[202:196];							
	assign ascii_6783_029 =ascii_IN[209:203];							
	assign ascii_6783_030 =ascii_IN[216:210];							
	assign ascii_6783_031 =ascii_IN[223:217];							
	assign ascii_6783_032 =ascii_IN[230:224];							
	assign ascii_6783_033 =ascii_IN[237:231];							
	assign ascii_6783_034 =ascii_IN[244:238];							
	assign ascii_6783_035 =ascii_IN[251:245];							
	assign ascii_6783_036 =ascii_IN[258:252];							
	assign ascii_6783_037 =ascii_IN[265:259];							
	assign ascii_6783_038 =ascii_IN[272:266];							
	assign ascii_6783_039 =ascii_IN[279:273];							
	assign ascii_6783_040 =ascii_IN[286:280];							
	assign ascii_6783_041 =ascii_IN[293:287];							
	assign ascii_6783_042 =ascii_IN[300:294];							
	assign ascii_6783_043 =ascii_IN[307:301];							
	assign ascii_6783_044 =ascii_IN[314:308];							
	assign ascii_6783_045 =ascii_IN[321:315];							
	assign ascii_6783_046 =ascii_IN[328:322];							
	assign ascii_6783_047 =ascii_IN[335:329];							
	assign ascii_6783_048 =ascii_IN[342:336];							
	assign ascii_6783_049 =ascii_IN[349:343];							
	assign ascii_6783_050 =ascii_IN[356:350];							
	assign ascii_6783_051 =ascii_IN[363:357];							
	assign ascii_6783_052 =ascii_IN[370:364];							
	assign ascii_6783_053 =ascii_IN[377:371];							
	assign ascii_6783_054 =ascii_IN[384:378];							
	assign ascii_6783_055 =ascii_IN[391:385];							
	assign ascii_6783_056 =ascii_IN[398:392];							
	assign ascii_6783_057 =ascii_IN[405:399];							
	assign ascii_6783_058 =ascii_IN[412:406];							
	assign ascii_6783_059 =ascii_IN[419:413];							
	assign ascii_6783_060 =ascii_IN[426:420];							
	assign ascii_6783_061 =ascii_IN[433:427];							
	assign ascii_6783_062 =ascii_IN[440:434];							
	assign ascii_6783_063 =ascii_IN[447:441];							
	assign ascii_6783_064 =ascii_IN[454:448];							
	assign ascii_6783_065 =ascii_IN[461:455];							
	assign ascii_6783_066 =ascii_IN[468:462];							
	assign ascii_6783_067 =ascii_IN[475:469];							
	assign ascii_6783_068 =ascii_IN[482:476];							
	assign ascii_6783_069 =ascii_IN[489:483];							
	assign ascii_6783_070 =ascii_IN[496:490];							
	assign ascii_6783_071 =ascii_IN[503:497];							
	assign ascii_6783_072 =ascii_IN[510:504];							
	assign ascii_6783_073 =ascii_IN[517:511];							
	assign ascii_6783_074 =ascii_IN[524:518];							
	assign ascii_6783_075 =ascii_IN[531:525];							
	assign ascii_6783_076 =ascii_IN[538:532];							
	assign ascii_6783_077 =ascii_IN[545:539];							
	assign ascii_6783_078 =ascii_IN[552:546];							
	assign ascii_6783_079 =ascii_IN[559:553];							
	assign ascii_6783_080 =ascii_IN[566:560];							
	assign ascii_6783_081 =ascii_IN[573:567];							
	assign ascii_6783_082 =ascii_IN[580:574];							
	assign ascii_6783_083 =ascii_IN[587:581];							
	assign ascii_6783_084 =ascii_IN[594:588];							
	assign ascii_6783_085 =ascii_IN[601:595];							
	assign ascii_6783_086 =ascii_IN[608:602];							
	assign ascii_6783_087 =ascii_IN[615:609];							
	assign ascii_6783_088 =ascii_IN[622:616];							
	assign ascii_6783_089 =ascii_IN[629:623];							
	assign ascii_6783_090 =ascii_IN[636:630];							
	assign ascii_6783_091 =ascii_IN[643:637];							

endmodule