module two_tgbase_to_one_big_number(
	input[5:0]	 tgBASE_6783_000,	tgBASE_6783_001,    tgBASE_6783_002,    tgBASE_6783_003,							
				 tgBASE_6783_004,	tgBASE_6783_005,	tgBASE_6783_006,	tgBASE_6783_007,	
				 tgBASE_6783_008,	tgBASE_6783_009,	tgBASE_6783_010,	tgBASE_6783_011,	
				 tgBASE_6783_012,	tgBASE_6783_013,	tgBASE_6783_014,	tgBASE_6783_015,	
				 tgBASE_6783_016,	tgBASE_6783_017,	tgBASE_6783_018,	tgBASE_6783_019,	
				 tgBASE_6783_020,	tgBASE_6783_021,	tgBASE_6783_022,	tgBASE_6783_023,	
				 tgBASE_6783_024,	tgBASE_6783_025,	tgBASE_6783_026,	tgBASE_6783_027,	
				 tgBASE_6783_028,	tgBASE_6783_029,	tgBASE_6783_030,	tgBASE_6783_031,	
				 tgBASE_6783_032,	tgBASE_6783_033,	tgBASE_6783_034,	tgBASE_6783_035,	
				 tgBASE_6783_036,	tgBASE_6783_037,	tgBASE_6783_038,	tgBASE_6783_039,	
				 tgBASE_6783_040,	tgBASE_6783_041,	tgBASE_6783_042,	tgBASE_6783_043,	
				 tgBASE_6783_044,	tgBASE_6783_045,	tgBASE_6783_046,	tgBASE_6783_047,	
				 tgBASE_6783_048,	tgBASE_6783_049,	tgBASE_6783_050,	tgBASE_6783_051,	
				 tgBASE_6783_052,	tgBASE_6783_053,	tgBASE_6783_054,	tgBASE_6783_055,	
				 tgBASE_6783_056,	tgBASE_6783_057,	tgBASE_6783_058,	tgBASE_6783_059,	
				 tgBASE_6783_060,	tgBASE_6783_061,	tgBASE_6783_062,	tgBASE_6783_063,	
				 tgBASE_6783_064,	tgBASE_6783_065,	tgBASE_6783_066,	tgBASE_6783_067,	
				 tgBASE_6783_068,	tgBASE_6783_069,	tgBASE_6783_070,	tgBASE_6783_071,	
				 tgBASE_6783_072,	tgBASE_6783_073,	tgBASE_6783_074,	tgBASE_6783_075,	
				 tgBASE_6783_076,	tgBASE_6783_077,	tgBASE_6783_078,	tgBASE_6783_079,	
				 tgBASE_6783_080,	tgBASE_6783_081,	tgBASE_6783_082,	tgBASE_6783_083,	
				 tgBASE_6783_084,	tgBASE_6783_085,	tgBASE_6783_086,	tgBASE_6783_087,	
				 tgBASE_6783_088,	tgBASE_6783_089,	tgBASE_6783_090,	tgBASE_6783_091,	
				 tgBASE_6783_092,	tgBASE_6783_093,	tgBASE_6783_094,	tgBASE_6783_095,	
				 tgBASE_6783_096,	tgBASE_6783_097,	tgBASE_6783_098,	tgBASE_6783_099,	
				 tgBASE_6783_100,	tgBASE_6783_101,	tgBASE_6783_102,	tgBASE_6783_103,	
				 tgBASE_6783_104,	tgBASE_6783_105,	tgBASE_6783_106,	tgBASE_6783_107,	
				 tgBASE_6783_108,	tgBASE_6783_109,	tgBASE_6783_110,	tgBASE_6783_111,	
				 tgBASE_6783_112,	tgBASE_6783_113,	tgBASE_6783_114,	tgBASE_6783_115,	
				 tgBASE_6783_116,	tgBASE_6783_117,	tgBASE_6783_118,	tgBASE_6783_119,	
				 tgBASE_6783_120,	tgBASE_6783_121,	tgBASE_6783_122,	tgBASE_6783_123,	
				 tgBASE_6783_124,	tgBASE_6783_125,	tgBASE_6783_126,	tgBASE_6783_127,	
				 tgBASE_6783_128,	tgBASE_6783_129,	tgBASE_6783_130,	tgBASE_6783_131,	
				 tgBASE_6783_132,	tgBASE_6783_133,	tgBASE_6783_134,	tgBASE_6783_135,	
				 tgBASE_6783_136,	tgBASE_6783_137,	tgBASE_6783_138,	tgBASE_6783_139,	
				 tgBASE_6783_140,	tgBASE_6783_141,	tgBASE_6783_142,	tgBASE_6783_143,	
				 tgBASE_6783_144,	tgBASE_6783_145,
	output[13:0] oneBig_6783_000,	oneBig_6783_001,    oneBig_6783_002,    oneBig_6783_003,							
				 oneBig_6783_004,	oneBig_6783_005,	oneBig_6783_006,	oneBig_6783_007,	
				 oneBig_6783_008,	oneBig_6783_009,	oneBig_6783_010,	oneBig_6783_011,	
				 oneBig_6783_012,	oneBig_6783_013,	oneBig_6783_014,	oneBig_6783_015,	
				 oneBig_6783_016,	oneBig_6783_017,	oneBig_6783_018,	oneBig_6783_019,	
				 oneBig_6783_020,	oneBig_6783_021,	oneBig_6783_022,	oneBig_6783_023,	
				 oneBig_6783_024,	oneBig_6783_025,	oneBig_6783_026,	oneBig_6783_027,	
				 oneBig_6783_028,	oneBig_6783_029,	oneBig_6783_030,	oneBig_6783_031,	
				 oneBig_6783_032,	oneBig_6783_033,	oneBig_6783_034,	oneBig_6783_035,	
				 oneBig_6783_036,	oneBig_6783_037,	oneBig_6783_038,	oneBig_6783_039,	
				 oneBig_6783_040,	oneBig_6783_041,	oneBig_6783_042,	oneBig_6783_043,	
				 oneBig_6783_044,	oneBig_6783_045,	oneBig_6783_046,	oneBig_6783_047,	
				 oneBig_6783_048,	oneBig_6783_049,	oneBig_6783_050,	oneBig_6783_051,	
				 oneBig_6783_052,	oneBig_6783_053,	oneBig_6783_054,	oneBig_6783_055,	
				 oneBig_6783_056,	oneBig_6783_057,	oneBig_6783_058,	oneBig_6783_059,	
				 oneBig_6783_060,	oneBig_6783_061,	oneBig_6783_062,	oneBig_6783_063,	
				 oneBig_6783_064,	oneBig_6783_065,	oneBig_6783_066,	oneBig_6783_067,	
				 oneBig_6783_068,	oneBig_6783_069,	oneBig_6783_070,	oneBig_6783_071,	
				 oneBig_6783_072);
				 
	assign oneBig_6783_000 =tgBASE_6783_000* 100 + tgBASE_6783_001;
	assign oneBig_6783_001 =tgBASE_6783_002* 100 + tgBASE_6783_003;
	assign oneBig_6783_002 =tgBASE_6783_004* 100 + tgBASE_6783_005;
	assign oneBig_6783_003 =tgBASE_6783_006* 100 + tgBASE_6783_007;
	assign oneBig_6783_004 =tgBASE_6783_008* 100 + tgBASE_6783_009;
	assign oneBig_6783_005 =tgBASE_6783_010* 100 + tgBASE_6783_011;
	assign oneBig_6783_006 =tgBASE_6783_012* 100 + tgBASE_6783_013;
	assign oneBig_6783_007 =tgBASE_6783_014* 100 + tgBASE_6783_015;
	assign oneBig_6783_008 =tgBASE_6783_016* 100 + tgBASE_6783_017;
	assign oneBig_6783_009 =tgBASE_6783_018* 100 + tgBASE_6783_019;
	assign oneBig_6783_010 =tgBASE_6783_020* 100 + tgBASE_6783_021;
	assign oneBig_6783_011 =tgBASE_6783_022* 100 + tgBASE_6783_023;
	assign oneBig_6783_012 =tgBASE_6783_024* 100 + tgBASE_6783_025;
	assign oneBig_6783_013 =tgBASE_6783_026* 100 + tgBASE_6783_027;
	assign oneBig_6783_014 =tgBASE_6783_028* 100 + tgBASE_6783_029;
	assign oneBig_6783_015 =tgBASE_6783_030* 100 + tgBASE_6783_031;
	assign oneBig_6783_016 =tgBASE_6783_032* 100 + tgBASE_6783_033;
	assign oneBig_6783_017 =tgBASE_6783_034* 100 + tgBASE_6783_035;
	assign oneBig_6783_018 =tgBASE_6783_036* 100 + tgBASE_6783_037;
	assign oneBig_6783_019 =tgBASE_6783_038* 100 + tgBASE_6783_039;
	assign oneBig_6783_020 =tgBASE_6783_040* 100 + tgBASE_6783_041;
	assign oneBig_6783_021 =tgBASE_6783_042* 100 + tgBASE_6783_043;
	assign oneBig_6783_022 =tgBASE_6783_044* 100 + tgBASE_6783_045;
	assign oneBig_6783_023 =tgBASE_6783_046* 100 + tgBASE_6783_047;
	assign oneBig_6783_024 =tgBASE_6783_048* 100 + tgBASE_6783_049;
	assign oneBig_6783_025 =tgBASE_6783_050* 100 + tgBASE_6783_051;
	assign oneBig_6783_026 =tgBASE_6783_052* 100 + tgBASE_6783_053;
	assign oneBig_6783_027 =tgBASE_6783_054* 100 + tgBASE_6783_055;
	assign oneBig_6783_028 =tgBASE_6783_056* 100 + tgBASE_6783_057;
	assign oneBig_6783_029 =tgBASE_6783_058* 100 + tgBASE_6783_059;
	assign oneBig_6783_030 =tgBASE_6783_060* 100 + tgBASE_6783_061;
	assign oneBig_6783_031 =tgBASE_6783_062* 100 + tgBASE_6783_063;
	assign oneBig_6783_032 =tgBASE_6783_064* 100 + tgBASE_6783_065;
	assign oneBig_6783_033 =tgBASE_6783_066* 100 + tgBASE_6783_067;
	assign oneBig_6783_034 =tgBASE_6783_068* 100 + tgBASE_6783_069;
	assign oneBig_6783_035 =tgBASE_6783_070* 100 + tgBASE_6783_071;
	assign oneBig_6783_036 =tgBASE_6783_072* 100 + tgBASE_6783_073;
	assign oneBig_6783_037 =tgBASE_6783_074* 100 + tgBASE_6783_075;
	assign oneBig_6783_038 =tgBASE_6783_076* 100 + tgBASE_6783_077;
	assign oneBig_6783_039 =tgBASE_6783_078* 100 + tgBASE_6783_079;
	assign oneBig_6783_040 =tgBASE_6783_080* 100 + tgBASE_6783_081;
	assign oneBig_6783_041 =tgBASE_6783_082* 100 + tgBASE_6783_083;
	assign oneBig_6783_042 =tgBASE_6783_084* 100 + tgBASE_6783_085;
	assign oneBig_6783_043 =tgBASE_6783_086* 100 + tgBASE_6783_087;
	assign oneBig_6783_044 =tgBASE_6783_088* 100 + tgBASE_6783_089;
	assign oneBig_6783_045 =tgBASE_6783_090* 100 + tgBASE_6783_091;
	assign oneBig_6783_046 =tgBASE_6783_092* 100 + tgBASE_6783_093;
	assign oneBig_6783_047 =tgBASE_6783_094* 100 + tgBASE_6783_095;
	assign oneBig_6783_048 =tgBASE_6783_096* 100 + tgBASE_6783_097;
	assign oneBig_6783_049 =tgBASE_6783_098* 100 + tgBASE_6783_099;
	assign oneBig_6783_050 =tgBASE_6783_100* 100 + tgBASE_6783_101;
	assign oneBig_6783_051 =tgBASE_6783_102* 100 + tgBASE_6783_103;
	assign oneBig_6783_052 =tgBASE_6783_104* 100 + tgBASE_6783_105;
	assign oneBig_6783_053 =tgBASE_6783_106* 100 + tgBASE_6783_107;
	assign oneBig_6783_054 =tgBASE_6783_108* 100 + tgBASE_6783_109;
	assign oneBig_6783_055 =tgBASE_6783_110* 100 + tgBASE_6783_111;
	assign oneBig_6783_056 =tgBASE_6783_112* 100 + tgBASE_6783_113;
	assign oneBig_6783_057 =tgBASE_6783_114* 100 + tgBASE_6783_115;
	assign oneBig_6783_058 =tgBASE_6783_116* 100 + tgBASE_6783_117;
	assign oneBig_6783_059 =tgBASE_6783_118* 100 + tgBASE_6783_119;
	assign oneBig_6783_060 =tgBASE_6783_120* 100 + tgBASE_6783_121;
	assign oneBig_6783_061 =tgBASE_6783_122* 100 + tgBASE_6783_123;
	assign oneBig_6783_062 =tgBASE_6783_124* 100 + tgBASE_6783_125;
	assign oneBig_6783_063 =tgBASE_6783_126* 100 + tgBASE_6783_127;
	assign oneBig_6783_064 =tgBASE_6783_128* 100 + tgBASE_6783_129;
	assign oneBig_6783_065 =tgBASE_6783_130* 100 + tgBASE_6783_131;
	assign oneBig_6783_066 =tgBASE_6783_132* 100 + tgBASE_6783_133;
	assign oneBig_6783_067 =tgBASE_6783_134* 100 + tgBASE_6783_135;
	assign oneBig_6783_068 =tgBASE_6783_136* 100 + tgBASE_6783_137;
	assign oneBig_6783_069 =tgBASE_6783_138* 100 + tgBASE_6783_139;
	assign oneBig_6783_070 =tgBASE_6783_140* 100 + tgBASE_6783_141;
	assign oneBig_6783_071 =tgBASE_6783_142* 100 + tgBASE_6783_143;
	assign oneBig_6783_072 =tgBASE_6783_144* 100 + tgBASE_6783_145;
endmodule